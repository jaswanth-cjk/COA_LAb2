`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:47:16 09/14/2022 
// Design Name: 
// Module Name:    B_4_bit_wrapper 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module B_4_bit_wrapper(input clk, input rst, output reg [3:0] y);



always @(posedge clk)
begin



end 

B_4_bit_upcounter ()
endmodule
